module keyboard_sim