module day(clk);
	input clk;





endmodule
