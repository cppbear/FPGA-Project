module show_count(mycount,seg5,seg6);
	input [7:0]mycount;
	output reg [6:0]seg5;
	output reg [6:0]seg6;
	
	always
	begin		
			case(mycount[3:0])
			0: seg5[6:0] = 7'b1000000;
			1: seg5[6:0] = 7'b1111001;
			2: seg5[6:0] = 7'b0100100;
			3: seg5[6:0] = 7'b0110000;
			4: seg5[6:0] = 7'b0011001;
			5: seg5[6:0] = 7'b0010010;
			6: seg5[6:0] = 7'b0000010;
			7: seg5[6:0] = 7'b1111000;
			8: seg5[6:0] = 7'b0000000;
			9: seg5[6:0] = 7'b0010000;
			10:seg5[6:0] = 7'b0001000;
			11:seg5[6:0] = 7'b0000011;
			12:seg5[6:0] = 7'b1000110;
			13:seg5[6:0] = 7'b0100001;
			14:seg5[6:0] = 7'b0000110;
			15:seg5[6:0] = 7'b0001110;
			default: seg5[6:0] = 7'b1000000;
			endcase
		
			case(mycount[7:4])
			0: seg6[6:0] = 7'b1000000;
			1: seg6[6:0] = 7'b1111001;
			2: seg6[6:0] = 7'b0100100;
			3: seg6[6:0] = 7'b0110000;
			4: seg6[6:0] = 7'b0011001;
			5: seg6[6:0] = 7'b0010010;
			6: seg6[6:0] = 7'b0000010;
			7: seg6[6:0] = 7'b1111000;
			8: seg6[6:0] = 7'b0000000;
			9: seg6[6:0] = 7'b0010000;
			10:seg6[6:0] = 7'b0001000;
			11:seg6[6:0] = 7'b0000011;
			12:seg6[6:0] = 7'b1000110;
			13:seg6[6:0] = 7'b0100001;
			14:seg6[6:0] = 7'b0000110;
			15:seg6[6:0] = 7'b0001110;
			default: seg6[6:0] = 7'b1000000;
			endcase
	end
endmodule

