module out_put(x, y1,y2,pre);
	input [7:0] x;
	output reg [6:0] y1;
	input pre;
	output reg [6:0] y2;
	always @(*)
	begin
		if(((pre == 1) && (x[7:0] != 8'hf0)))	
		begin	
			case(x[3:0])
			0: y1[6:0] = 7'b1000000;
			1: y1[6:0] = 7'b1111001;
			2: y1[6:0] = 7'b0100100;
			3: y1[6:0] = 7'b0110000;
			4: y1[6:0] = 7'b0011001;
			5: y1[6:0] = 7'b0010010;
			6: y1[6:0] = 7'b0000010;
			7: y1[6:0] = 7'b1111000;
			8: y1[6:0] = 7'b0000000;
			9: y1[6:0] = 7'b0010000;
			10:y1[6:0] = 7'b0001000;
			11:y1[6:0] = 7'b0000011;
			12:y1[6:0] = 7'b1000110;
			13:y1[6:0] = 7'b0100001;
			14:y1[6:0] = 7'b0000110;
			15:y1[6:0] = 7'b0001110;
			endcase
		
			case(x[7:4])
			0: y2[6:0] = 7'b1000000;
			1: y2[6:0] = 7'b1111001;
			2: y2[6:0] = 7'b0100100;
			3: y2[6:0] = 7'b0110000;
			4: y2[6:0] = 7'b0011001;
			5: y2[6:0] = 7'b0010010;
			6: y2[6:0] = 7'b0000010;
			7: y2[6:0] = 7'b1111000;
			8: y2[6:0] = 7'b0000000;
			9: y2[6:0] = 7'b0010000;
			10:y2[6:0] = 7'b0001000;
			11:y2[6:0] = 7'b0000011;
			12:y2[6:0] = 7'b1000110;
			13:y2[6:0] = 7'b0100001;
			14:y2[6:0] = 7'b0000110;
			15:y2[6:0] = 7'b0001110;
			endcase
		end
		else
		begin
			y1[6:0] = 7'b1111111;
			y2[6:0] = 7'b1111111;
		end
	end
	
endmodule 