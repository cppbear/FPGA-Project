module picture(clk, reset, clken, vga_clk, hsync, vsync, valid, red, green, blue);
	input clk, reset, clken;
	reg [23:0] data=24'b0;
	output vga_clk, hsync, vsync, valid;
	wire temp_clk;
	wire [9:0] h_addr, v_addr;
	output [7:0] red, green, blue;
	reg [18:0] rom_addr=19'b0;
	wire [11:0] temp_color;
	
	clkgen #(25000000) clk_(clk, 1'b0, 1'b1, temp_clk);
	vga_ctrl ctrl(temp_clk, 1'b0, data, h_addr, v_addr, hsync, vsync, valid, red, green, blue);
	ROM rom(rom_addr, temp_clk, temp_color);
	assign vga_clk = temp_clk;
	
	always @(posedge clk)
	begin
		rom_addr = {h_addr, v_addr[8:0]};
		data[23:20] = temp_color[11:8];
		data[19:16] = 4'b0000;
		data[15:12] = temp_color[7:4];
		data[11:8] = 4'b0000;
		data[7:4] = temp_color[3:0];
		data[3:0] = 4'b0000;
	end

endmodule
