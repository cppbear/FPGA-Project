module show (pre,my_data,seg1,seg2,preflag);
	input pre;
	input preflag;
	input [7:0] my_data;
	output reg [6:0]seg1;
	output reg [6:0]seg2;
	
	always
	begin
		if(((pre == 1) && (my_data[7:0] != 8'hf0)))	
		begin	
			case(my_data[3:0])
			0: seg1[6:0] = 7'b1000000;
			1: seg1[6:0] = 7'b1111001;
			2: seg1[6:0] = 7'b0100100;
			3: seg1[6:0] = 7'b0110000;
			4: seg1[6:0] = 7'b0011001;
			5: seg1[6:0] = 7'b0010010;
			6: seg1[6:0] = 7'b0000010;
			7: seg1[6:0] = 7'b1111000;
			8: seg1[6:0] = 7'b0000000;
			9: seg1[6:0] = 7'b0010000;
			10:seg1[6:0] = 7'b0001000;
			11:seg1[6:0] = 7'b0000011;
			12:seg1[6:0] = 7'b1000110;
			13:seg1[6:0] = 7'b0100001;
			14:seg1[6:0] = 7'b0000110;
			15:seg1[6:0] = 7'b0001110;
			endcase
		
			case(my_data[7:4])
			0: seg2[6:0] = 7'b1000000;
			1: seg2[6:0] = 7'b1111001;
			2: seg2[6:0] = 7'b0100100;
			3: seg2[6:0] = 7'b0110000;
			4: seg2[6:0] = 7'b0011001;
			5: seg2[6:0] = 7'b0010010;
			6: seg2[6:0] = 7'b0000010;
			7: seg2[6:0] = 7'b1111000;
			8: seg2[6:0] = 7'b0000000;
			9: seg2[6:0] = 7'b0010000;
			10:seg2[6:0] = 7'b0001000;
			11:seg2[6:0] = 7'b0000011;
			12:seg2[6:0] = 7'b1000110;
			13:seg2[6:0] = 7'b0100001;
			14:seg2[6:0] = 7'b0000110;
			15:seg2[6:0] = 7'b0001110;
			endcase
		end
		else
		begin
			seg1[6:0] = 7'b1111111;
			seg2[6:0] = 7'b1111111;
		end
	end
endmodule
